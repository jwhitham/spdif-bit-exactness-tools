
library ieee;
use ieee.std_logic_1164.all;

entity test_signal_generator is
    port (
        data        : out std_logic
    );
end test_signal_generator;

architecture structural of test_signal_generator is
begin
    process
    begin
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '0';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '1';
wait for 80 ns;
data <= '0';

        wait;
    end;
end structural;
