
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity match_rom is
    port (
        address_in       : in std_logic_vector (6 downto 0) := (others => '0');
        data_out         : out std_logic_vector (23 downto 0) := (others => '0');
        clock            : in std_logic
    );
end match_rom;

architecture structural of match_rom is
begin
    process (clock)
    begin
        if clock = '1' and clock'event then
            case address_in is
when "0000000" => data_out <= "000000000000000000000000";
when "0000001" => data_out <= "011001010100001100100001";
when "0000010" => data_out <= "110001100100111000000000";
when "0000011" => data_out <= "011001010101111000000000";
when "0000100" => data_out <= "001001010111011000000000";
when "0000101" => data_out <= "011111010101011000000000";
when "0000110" => data_out <= "111101100110100100000000";
when "0000111" => data_out <= "010100011111001100000000";
when "0001000" => data_out <= "101101100001100000000000";
when "0001001" => data_out <= "000111010111011000000000";
when "0001010" => data_out <= "010011011100000100000000";
when "0001011" => data_out <= "110110110101111000000000";
when "0001100" => data_out <= "010000001101100100000000";
when "0001101" => data_out <= "100111100000110100000000";
when "0001110" => data_out <= "010100001000101000000000";
when "0001111" => data_out <= "010010001101110100000000";
when "0010000" => data_out <= "111000111011001100001101";
when "0010001" => data_out <= "000011001000111110101111";
when "0010010" => data_out <= "101011111110011001011110";
when "0010011" => data_out <= "010000011001010110110011";
when "0010100" => data_out <= "011001100111000000000001";
when "0010101" => data_out <= "010000001000000101111111";
when "0010110" => data_out <= "001001001101101011110001";
when "0010111" => data_out <= "111010111111100011001001";
when "0011000" => data_out <= "010110100010000011001001";
when "0011001" => data_out <= "011101011100001111101010";
when "0011010" => data_out <= "110100001001011000011100";
when "0011011" => data_out <= "100011011110001110110011";
when "0011100" => data_out <= "100011111011010000001000";
when "0011101" => data_out <= "110011111011010101010101";
when "0011110" => data_out <= "111010100110110101100110";
when "0011111" => data_out <= "001111100100100001110100";
when "0100000" => data_out <= "000000000000000000000001";
when "0100001" => data_out <= "111111111111111111111110";
when "0100010" => data_out <= "000000000000000000000010";
when "0100011" => data_out <= "111111111111111111111101";
when "0100100" => data_out <= "000000000000000000000100";
when "0100101" => data_out <= "111111111111111111111011";
when "0100110" => data_out <= "000000000000000000001000";
when "0100111" => data_out <= "111111111111111111110111";
when "0101000" => data_out <= "000000000000000000010000";
when "0101001" => data_out <= "111111111111111111101111";
when "0101010" => data_out <= "000000000000000000100000";
when "0101011" => data_out <= "111111111111111111011111";
when "0101100" => data_out <= "000000000000000001000000";
when "0101101" => data_out <= "111111111111111110111111";
when "0101110" => data_out <= "000000000000000010000000";
when "0101111" => data_out <= "111111111111111101111111";
when "0110000" => data_out <= "000000000000000100000000";
when "0110001" => data_out <= "111111111111111011111111";
when "0110010" => data_out <= "000000000000001000000000";
when "0110011" => data_out <= "111111111111110111111111";
when "0110100" => data_out <= "000000000000010000000000";
when "0110101" => data_out <= "111111111111101111111111";
when "0110110" => data_out <= "000000000000100000000000";
when "0110111" => data_out <= "111111111111011111111111";
when "0111000" => data_out <= "000000000001000000000000";
when "0111001" => data_out <= "111111111110111111111111";
when "0111010" => data_out <= "000000000010000000000000";
when "0111011" => data_out <= "111111111101111111111111";
when "0111100" => data_out <= "000000000100000000000000";
when "0111101" => data_out <= "111111111011111111111111";
when "0111110" => data_out <= "000000001000000000000000";
when "0111111" => data_out <= "111111110111111111111111";
when "1000000" => data_out <= "000000010000000000000000";
when "1000001" => data_out <= "111111101111111111111111";
when "1000010" => data_out <= "000000100000000000000000";
when "1000011" => data_out <= "111111011111111111111111";
when "1000100" => data_out <= "000001000000000000000000";
when "1000101" => data_out <= "111110111111111111111111";
when "1000110" => data_out <= "000010000000000000000000";
when "1000111" => data_out <= "111101111111111111111111";
when "1001000" => data_out <= "000100000000000000000000";
when "1001001" => data_out <= "111011111111111111111111";
when "1001010" => data_out <= "001000000000000000000000";
when "1001011" => data_out <= "110111111111111111111111";
when "1001100" => data_out <= "010000000000000000000000";
when "1001101" => data_out <= "101111111111111111111111";
when "1001110" => data_out <= "100000000000000000000000";
when "1001111" => data_out <= "011111111111111111111111";
when others =>   data_out <= "000000000000000000000000";

            end case;
        end if;
    end process;
end structural;
