package filter_unit_settings is
constant FRACTIONAL_BITS : Natural := 14;
constant NON_FRACTIONAL_BITS : Natural := 2;
constant UC_ADDR_BITS : Natural := 9;
constant ALL_BITS : Natural := 16;
constant A_BITS : Natural := 30;
constant VERBOSE_DEBUG : Boolean := False;
constant DATA_BITS : Natural := 16;
constant BAUD_RATE : Real := 300.0;
constant SAMPLE_RATE : Real := 48000.0;

end package filter_unit_settings;
