
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity filter_unit_microcode_store is port (
        uc_data_out : out std_logic_vector (7 downto 0) := (others => '0');
        uc_addr_in  : in std_logic_vector (8 downto 0) := (others => '0');
        enable_in   : in std_logic := '0';
        clock_in    : in std_logic := '0');
end filter_unit_microcode_store;
architecture behavioural of filter_unit_microcode_store is
    subtype t_word is std_logic_vector (7 downto 0);
    type t_storage is array (0 to 511) of t_word;
    signal storage : t_storage := (
0 => "00000001",
1 => "11000100",
2 => "10000000",
3 => "01100000",
4 => "10000111",
5 => "11000010",
6 => "00100010",
7 => "00100010",
8 => "00100010",
9 => "00100010",
10 => "00100010",
11 => "00100010",
12 => "00100010",
13 => "00100010",
14 => "00100010",
15 => "00100010",
16 => "00100010",
17 => "00100010",
18 => "00100010",
19 => "00100010",
20 => "00100010",
21 => "00100000",
22 => "00100000",
23 => "00100000",
24 => "00100000",
25 => "00100000",
26 => "00100000",
27 => "00100000",
28 => "00100000",
29 => "00100000",
30 => "00100011",
31 => "00100011",
32 => "00100000",
33 => "00100000",
34 => "00100000",
35 => "00100000",
36 => "00100010",
37 => "10000000",
38 => "01100000",
39 => "01100000",
40 => "11000011",
41 => "10001001",
42 => "11000010",
43 => "00100100",
44 => "00100101",
45 => "00100101",
46 => "00100101",
47 => "00100101",
48 => "00100101",
49 => "00100101",
50 => "00100101",
51 => "00100101",
52 => "00100101",
53 => "00100101",
54 => "00100101",
55 => "00100101",
56 => "00100101",
57 => "00100101",
58 => "00100011",
59 => "00100011",
60 => "00100011",
61 => "00100011",
62 => "00100011",
63 => "00100011",
64 => "00100011",
65 => "00100011",
66 => "00100011",
67 => "00100000",
68 => "00100011",
69 => "00100000",
70 => "00100000",
71 => "00100000",
72 => "00100000",
73 => "00100100",
74 => "10000000",
75 => "01100000",
76 => "01100000",
77 => "11000011",
78 => "10000011",
79 => "11000010",
80 => "00100110",
81 => "00100111",
82 => "00100111",
83 => "00100111",
84 => "00100111",
85 => "00100111",
86 => "00100111",
87 => "00100111",
88 => "00100111",
89 => "00100111",
90 => "00100111",
91 => "00100111",
92 => "00100111",
93 => "00100111",
94 => "00100111",
95 => "00100011",
96 => "00100000",
97 => "00100000",
98 => "00100000",
99 => "00100000",
100 => "00100011",
101 => "00100000",
102 => "00100011",
103 => "00100000",
104 => "00100000",
105 => "00100000",
106 => "00100011",
107 => "00100000",
108 => "00100011",
109 => "00100011",
110 => "00100110",
111 => "10000000",
112 => "01100000",
113 => "01100000",
114 => "11000011",
115 => "10000100",
116 => "11000010",
117 => "00101000",
118 => "00101001",
119 => "00101001",
120 => "00101001",
121 => "00101001",
122 => "00101001",
123 => "00101001",
124 => "00101001",
125 => "00101001",
126 => "00101001",
127 => "00101001",
128 => "00101001",
129 => "00101001",
130 => "00101001",
131 => "00101001",
132 => "00100011",
133 => "00100011",
134 => "00100000",
135 => "00100000",
136 => "00100000",
137 => "00100000",
138 => "00100000",
139 => "00100000",
140 => "00100011",
141 => "00100011",
142 => "00100000",
143 => "00100000",
144 => "00100000",
145 => "00100000",
146 => "00100000",
147 => "00101000",
148 => "10000011",
149 => "01001010",
150 => "00001011",
151 => "00001011",
152 => "00001011",
153 => "00001011",
154 => "00001011",
155 => "00001011",
156 => "00001011",
157 => "00001011",
158 => "00001011",
159 => "00001011",
160 => "00001011",
161 => "00001011",
162 => "00001011",
163 => "00001011",
164 => "10000001",
165 => "01001100",
166 => "11000100",
167 => "11000100",
168 => "10000000",
169 => "01100000",
170 => "10000110",
171 => "11000010",
172 => "00101101",
173 => "00101101",
174 => "00101101",
175 => "00101101",
176 => "00101101",
177 => "00101101",
178 => "00101101",
179 => "00101101",
180 => "00101101",
181 => "00101101",
182 => "00101101",
183 => "00101101",
184 => "00101101",
185 => "00101101",
186 => "00101101",
187 => "00100000",
188 => "00100000",
189 => "00100011",
190 => "00100011",
191 => "00100011",
192 => "00100011",
193 => "00100011",
194 => "00100011",
195 => "00100000",
196 => "00100000",
197 => "00100000",
198 => "00100011",
199 => "00100000",
200 => "00100011",
201 => "00100011",
202 => "00101101",
203 => "00001011",
204 => "00001011",
205 => "00001011",
206 => "00001011",
207 => "00001011",
208 => "00001011",
209 => "00001011",
210 => "00001011",
211 => "00001011",
212 => "00001011",
213 => "00001011",
214 => "00001011",
215 => "00001011",
216 => "00001011",
217 => "10000001",
218 => "01001110",
219 => "11000100",
220 => "11000100",
221 => "10000011",
222 => "00001111",
223 => "01010000",
224 => "11000001",
225 => "10000110",
226 => "00010001",
227 => "01010010",
228 => "11000001",
229 => "11000101",
230 => "10001111",
231 => "00010001",
232 => "01010011",
233 => "11000001",
234 => "11000100",
235 => "11000110",
236 => "11000111",
237 => "10001110",
238 => "11000100",
239 => "10000000",
240 => "01100000",
241 => "10000111",
242 => "11000010",
243 => "00100010",
244 => "00100010",
245 => "00100010",
246 => "00100010",
247 => "00100010",
248 => "00100010",
249 => "00100010",
250 => "00100010",
251 => "00100010",
252 => "00100010",
253 => "00100010",
254 => "00100010",
255 => "00100010",
256 => "00100010",
257 => "00100010",
258 => "00100000",
259 => "00100000",
260 => "00100000",
261 => "00100000",
262 => "00100000",
263 => "00100000",
264 => "00100000",
265 => "00100000",
266 => "00100011",
267 => "00100000",
268 => "00100000",
269 => "00100011",
270 => "00100000",
271 => "00100011",
272 => "00100000",
273 => "00100010",
274 => "10000000",
275 => "01100000",
276 => "01100000",
277 => "11000011",
278 => "10001001",
279 => "11000010",
280 => "00100100",
281 => "00100101",
282 => "00100101",
283 => "00100101",
284 => "00100101",
285 => "00100101",
286 => "00100101",
287 => "00100101",
288 => "00100101",
289 => "00100101",
290 => "00100101",
291 => "00100101",
292 => "00100101",
293 => "00100101",
294 => "00100101",
295 => "00100011",
296 => "00100011",
297 => "00100011",
298 => "00100011",
299 => "00100011",
300 => "00100011",
301 => "00100011",
302 => "00100011",
303 => "00100000",
304 => "00100011",
305 => "00100011",
306 => "00100000",
307 => "00100011",
308 => "00100011",
309 => "00100000",
310 => "00100100",
311 => "10000000",
312 => "01100000",
313 => "01100000",
314 => "11000011",
315 => "10000011",
316 => "11000010",
317 => "00100110",
318 => "00100111",
319 => "00100111",
320 => "00100111",
321 => "00100111",
322 => "00100111",
323 => "00100111",
324 => "00100111",
325 => "00100111",
326 => "00100111",
327 => "00100111",
328 => "00100111",
329 => "00100111",
330 => "00100111",
331 => "00100111",
332 => "00100011",
333 => "00100000",
334 => "00100000",
335 => "00100000",
336 => "00100011",
337 => "00100000",
338 => "00100011",
339 => "00100000",
340 => "00100011",
341 => "00100011",
342 => "00100000",
343 => "00100011",
344 => "00100000",
345 => "00100000",
346 => "00100000",
347 => "00100110",
348 => "10000000",
349 => "01100000",
350 => "01100000",
351 => "11000011",
352 => "10000100",
353 => "11000010",
354 => "00101000",
355 => "00101001",
356 => "00101001",
357 => "00101001",
358 => "00101001",
359 => "00101001",
360 => "00101001",
361 => "00101001",
362 => "00101001",
363 => "00101001",
364 => "00101001",
365 => "00101001",
366 => "00101001",
367 => "00101001",
368 => "00101001",
369 => "00100011",
370 => "00100011",
371 => "00100000",
372 => "00100000",
373 => "00100000",
374 => "00100000",
375 => "00100000",
376 => "00100011",
377 => "00100000",
378 => "00100000",
379 => "00100011",
380 => "00100000",
381 => "00100011",
382 => "00100000",
383 => "00100000",
384 => "00101000",
385 => "10000011",
386 => "01001010",
387 => "00001011",
388 => "00001011",
389 => "00001011",
390 => "00001011",
391 => "00001011",
392 => "00001011",
393 => "00001011",
394 => "00001011",
395 => "00001011",
396 => "00001011",
397 => "00001011",
398 => "00001011",
399 => "00001011",
400 => "00001011",
401 => "10000001",
402 => "01001100",
403 => "11000100",
404 => "11000100",
405 => "10000000",
406 => "01100000",
407 => "10000110",
408 => "11000010",
409 => "00101101",
410 => "00101101",
411 => "00101101",
412 => "00101101",
413 => "00101101",
414 => "00101101",
415 => "00101101",
416 => "00101101",
417 => "00101101",
418 => "00101101",
419 => "00101101",
420 => "00101101",
421 => "00101101",
422 => "00101101",
423 => "00101101",
424 => "00100000",
425 => "00100000",
426 => "00100011",
427 => "00100011",
428 => "00100011",
429 => "00100011",
430 => "00100011",
431 => "00100011",
432 => "00100000",
433 => "00100000",
434 => "00100000",
435 => "00100011",
436 => "00100000",
437 => "00100011",
438 => "00100011",
439 => "00101101",
440 => "00001011",
441 => "00001011",
442 => "00001011",
443 => "00001011",
444 => "00001011",
445 => "00001011",
446 => "00001011",
447 => "00001011",
448 => "00001011",
449 => "00001011",
450 => "00001011",
451 => "00001011",
452 => "00001011",
453 => "00001011",
454 => "10000001",
455 => "01001110",
456 => "11000100",
457 => "11000100",
458 => "10000011",
459 => "00001111",
460 => "01010000",
461 => "11000001",
462 => "10000110",
463 => "00010001",
464 => "01010010",
465 => "11000001",
466 => "11000101",
467 => "10001111",
468 => "00010001",
469 => "01010011",
470 => "11000001",
471 => "11000100",
472 => "11000110",
473 => "11000111",
474 => "10000110",
475 => "00010100",
476 => "01010011",
477 => "10001110",
478 => "10000110",
479 => "00010001",
480 => "01010010",
481 => "11000101",
482 => "00010101",
483 => "10001000",
484 => "01010110",
485 => "10000111",
486 => "01010111",
487 => "00011000",
others => x"ff");

begin
    process (clock_in)
    begin
        if clock_in'event and clock_in = '1' then
            if enable_in = '1' then
                uc_data_out <= storage (to_integer (unsigned (uc_addr_in)));
            end if;
        end if;
    end process;
end architecture behavioural;
