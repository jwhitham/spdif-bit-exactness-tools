spdif_out_pll_inst: spdif_out_pll
port map(
          REFERENCECLK => ,
          PLLOUTCORE => ,
          PLLOUTGLOBAL => ,
          RESET => ,
          LOCK => 
        );
