spdif_meter_pll_inst: spdif_meter_pll
port map(
          REFERENCECLK => ,
          PLLOUTCORE => ,
          PLLOUTGLOBAL => ,
          RESET => 
        );
